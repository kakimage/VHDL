entity is