library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
 
ENTITY ACC_TB IS
END ACC_TB;
 
ARCHITECTURE Behavioral OF ACC_TB IS
 
 COMPONENT ACC
 PORT(
		i_CLK : IN STD_LOGIC; 			
		i_RST : IN STD_LOGIC;
		i_WR_ACC : IN STD_LOGIC;
		i_ACC : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
		o_ACC : OUT STD_LOGIC_VECTOR (15 DOWNTO 0)
 );
 END COMPONENT;
 
 SIGNAL w_CLK : STD_LOGIC := '0';
 SIGNAL w_RST : STD_LOGIC := '0';
 SIGNAL w_WR_ACC: STD_LOGIC;
 SIGNAL wi_ACC : STD_LOGIC_VECTOR(15 downto 0) := (others => '0');
 
 SIGNAL wo_ACC : std_logic_vector(15 downto 0);
 
 
BEGIN
 
	UUT: ACC 
		PORT MAP (
		 i_CLK => w_CLK,
		 i_RST => w_RST,
		 i_WR_ACC => w_WR_ACC,
		 i_ACC => wi_ACC,
		 o_ACC => wo_ACC
		);

	--PROCESSO DE RELOGIO
	PROCESS
	BEGIN
		 w_CLK <= '0';
		 WAIT FOR 20 ns;
		 w_CLK <= '1';
		 WAIT FOR 20 ns;
	END PROCESS;
	 
	--CIRCUITO DE RESET 
	PROCESS
	BEGIN
		w_RST <= '1';
		WAIT FOR 100 ns;
		w_RST <= '0';
		WAIT;

	END PROCESS;
	
	--TESTE ACC
	PROCESS
	BEGIN
		wi_ACC <= "0000000000000001";
		WAIT FOR 150 ns;
		w_WR_ACC <= '1';
		WAIT;
	END PROCESS;
 
END Behavioral;
