library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


entity SETE_SEGMENTOS is
	 Port ( 
				i_NUMERO		: in  STD_LOGIC_VECTOR(3 DOWNTO 0);
				i_RST 		: in  STD_LOGIC;
			   o_DISPLAY  	: out STD_LOGIC_VECTOR(6 DOWNTO 0)
	 );
end SETE_SEGMENTOS;


architecture Behavioral of SETE_SEGMENTOS is


begin


	
end Behavioral;