LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
  
ENTITY TB_ULA IS
END TB_ULA;
  
ARCHITECTURE behavior OF TB_ULA IS
  
	COMPONENT ULA is
	PORT(
		i_INPUT_A : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		i_INPUT_B : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		i_INPUT_IR: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		i_SEL : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		o_OUTPUT : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
	END COMPONENT;
  
 
 signal i_INPUT_A : STD_LOGIC_VECTOR(15 DOWNTO 0) := (others => '0');
 signal i_INPUT_B : STD_LOGIC_VECTOR(3 DOWNTO 0) := (others => '0');
 signal i_INPUT_IR : STD_LOGIC_VECTOR(3 DOWNTO 0) := (others => '0');
 signal i_SEL : STD_LOGIC_VECTOR(2 DOWNTO 0) := (others => '0');
 
 signal o_OUTPUT : STD_LOGIC_VECTOR(15 DOWNTO 0);
  
BEGIN
  
	UUT: ULA PORT MAP (
		i_INPUT_A => i_INPUT_A,
		i_INPUT_B => i_INPUT_B,
		i_INPUT_IR => i_INPUT_IR,
		o_OUTPUT => o_OUTPUT
	);

	PROCESS
	BEGIN
	
	WAIT FOR 100 ns;

	i_INPUT_A <= "0000111100001001";
	i_INPUT_B <= "0000111100001111";
	i_INPUT_IR <= "0000111100001100";

	i_SEL <= "100";
	WAIT FOR 100 ns;
	i_SEL <= "101";
	WAIT FOR 100 ns;
	i_SEL <= "110";
	WAIT FOR 100 ns;
	i_SEL <= "111";

	end process;
 
END;
