library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use iEEE.NUMERIC_STD.ALL;

entity CONTROL is
	port(
		i_OPCODE: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		o_WR_RAM: OUT STD_LOGIC;
		o_EN_RAM: OUT STD_LOGIC;
		o_EN_PC: OUT STD_LOGIC;
		o_EN_ROM: OUT STD_LOGIC;
		o_WR_ACC: OUT STD_LOGIC;
		o_SEL_OP1: OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
		o_SEL_OP2: OUT STD_LOGIC;
		o_SEL_ULA: OUT STD_LOGIC;
		o_EN_IN: OUT STD_LOGIC
	);
end CONTROL;

architecture Behavioral of CONTROL is
	SIGNAL w_WR_RAM: STD_LOGIC;
	SIGNAL w_EN_RAM: STD_LOGIC;
	SIGNAL w_EN_PC: STD_LOGIC;
	SIGNAL w_EN_ROM: STD_LOGIC;
	SIGNAL w_WR_ACC: STD_LOGIC;
	SIGNAL w_SEL_OP1: STD_LOGIC_VECTOR(1 DOWNTO 0);
	SIGNAL w_SEL_OP2: STD_LOGIC;
	SIGNAL w_SEL_ULA: STD_LOGIC;
	SIGNAL w_EN_IN: STD_LOGIC;
	
begin
	w_WR_RAM <= (NOT i_OPCODE(3) AND NOT i_OPCODE(2) AND NOT i_OPCODE(1) AND i_OPCODE(0));
	w_EN_RAM <= ((NOT i_OPCODE(3) AND (NOT i_OPCODE(2) AND (i_OPCODE(1) XOR i_OPCODE(0)))) OR (i_OPCODE(2) AND NOT i_OPCODE(0)));
	w_EN_PC <= (i_OPCODE(3) OR i_OPCODE(2) or i_OPCODE(1) or i_OPCODE(0));
	w_EN_ROM <= w_EN_PC;
	w_WR_ACC <= (i_OPCODE(3) OR i_OPCODE(2) OR i_OPCODE(1));
	w_SEL_OP1(1) <= ((NOT i_OPCODE(3) AND i_OPCODE(2)) OR (i_OPCODE(3) AND NOT i_OPCODE(2) AND NOT i_OPCODE(1) AND i_OPCODE(0)));
	w_SEL_OP1(0) <= (NOT i_OPCODE(2) AND i_OPCODE(0));
	w_SEL_OP2 <= ((NOT i_OPCODE(2) AND i_OPCODE(0)) OR (NOT i_OPCODE(3) AND i_OPCODE(2) AND i_OPCODE(0)));
	w_SEL_ULA <= (NOT i_OPCODE(3) AND i_OPCODE(2) AND i_OPCODE(1));
	w_EN_IN <= (NOT i_OPCODE(3) AND i_OPCODE(2) AND i_OPCODE(1) AND NOT i_OPCODE(0));
	
	o_WR_RAM <= w_WR_RAM;
	o_EN_RAM <= w_EN_RAM;
	o_EN_PC <= w_EN_PC;
	o_EN_ROM <= w_EN_ROM;
	o_WR_ACC <= w_WR_ACC;
	o_SEL_OP1 <= w_SEL_OP1;
	o_SEL_OP2 <= w_SEL_OP2;
	o_SEL_ULA <= w_SEL_ULA;
	o_EN_IN <= w_EN_IN;
	
end Behavioral;