MULTIPLEX_inst : MULTIPLEX PORT MAP (
		clock	 => clock_sig,
		data_in	 => data_in_sig,
		sload_data	 => sload_data_sig,
		result	 => result_sig,
		result_valid	 => result_valid_sig
	);
