LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY FULL_ADDER IS
	PORT(
		I_A : IN  STD_LOGIC;
		I_B : IN  STD_LOGIC;
		I_C : IN  STD_LOGIC;
		O_C : OUT STD_LOGIC;
		O_S : OUT STD_LOGIC
	);
END ENTITY;

ARCHITECTURE BEHAVIORAL OF FULL_ADDER IS
	COMPONENT HALF_ADDER IS
		PORT(
			I_A : IN  STD_LOGIC;
			I_B : IN  STD_LOGIC;
			O_C : OUT STD_LOGIC;
			O_S : OUT STD_LOGIC
		);
	END COMPONENT;

	SIGNAL W_C1 : STD_LOGIC;
	SIGNAL W_C2 : STD_LOGIC;
	SIGNAL W_s  : STD_LOGIC;
BEGIN
	HALF1 : HALF_ADDER
	PORT MAP (
		I_A	=> I_A,
		I_B	=> I_B,
		O_S	=> W_S,
		O_C	=> W_C1
	);

	HALF2 : HALF_ADDER
	PORT MAP (
		I_A	=> W_S,
		I_B	=> I_C,
		O_S	=> O_S,
		O_C	=> W_C2
	);

	O_C <= W_C1 OR W_C2;
END ARCHITECTURE;