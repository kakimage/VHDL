LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY HALF_ADDER IS
	PORT(
        I_A : IN  STD_LOGIC;
        I_B : IN  STD_LOGIC;
        O_C : OUT STD_LOGIC;
        O_S : OUT STD_LOGIC
	);
END ENTITY;

ARCHITECTURE BEHAVIORAL OF HALF_ADDER IS

BEGIN
    O_S <= I_A XOR I_B;
    O_C <= I_A AND I_B;
END ARCHITECTURE;